module ex2(
	input [7:0]in,
	input en,
	output reg [2:0]out,
	output reg [6:0]out_hex0
);
	always@(*) begin
  		if (en) begin
  			casez (in)
  				8'b1???????: out = 3'b111;
        			8'b01??????: out = 3'b110;
        			8'b001?????: out = 3'b101;
        			8'b0001????: out = 3'b100;
        			8'b00001???: out = 3'b011;
        			8'b000001??: out = 3'b010;
        			8'b0000001?: out = 3'b001;
        			8'b00000001: out = 3'b000;
        			default:     out = 3'b000;
        		endcase
		end
		else begin
			out = 3'b000;
		end
		if(en) begin
			case(out)
				3'b111: out_hex0 = 7'b1111000;
				3'b110: out_hex0 = 7'b0000010;
				3'b101: out_hex0 = 7'b0001010;
				3'b100: out_hex0 = 7'b0011001;
				3'b011: out_hex0 = 7'b0110000;
				3'b010: out_hex0 = 7'b0100100;
				3'b001: out_hex0 = 7'b1111001;
				3'b000: out_hex0 = 7'b1000000;
				default:out_hex0 = 7'b1000000;
			endcase
		end
	end
endmodule
